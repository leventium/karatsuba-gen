module karatsuba_leaf_2x2 (
  input  [1:0] u, v,

  output [3:0] r
);

  assign r = u * v;

endmodule
